module next_state_gen(
    input x,
    input [1:0] q,
    output [1:0] x
)