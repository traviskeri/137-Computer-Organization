`include "multi_cycle_circuit.v"

module tester();

reg clock, reset, a, b, c, d;